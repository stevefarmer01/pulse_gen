package pulse_generator_pkg;

  const int blah = 0;

  localparam  reset_delay_c = 4;
  localparam  start_delay_c = 4;
  localparam  pulse_width_c = 4;

endpackage
